module Traffic_Light_Control_2 (
input wire clk, rs,
output reg [2:0] out_1, out_2
);

reg [1:0] Current_State, Next_State;
reg [4:0] t;
parameter S0 = 0, S1 = 1, S2 = 2, S3 = 3;
parameter Time_S0 = 15, Time_S1 = 5, Time_S2 = 15, Time_S3 = 5;

always @(posedge clk) begin
	if (rs) begin
		t <= Time_S0;
	end else if (t == 0) begin
		case (Next_State)
		S0: t <= Time_S0;
		S1: t <= Time_S1;
		S2: t <= Time_S2;
		S3: t <= Time_S3;
		default: t <= Time_S0;
	endcase
	end else begin
		t <= t - 1;
	end
end

always @(posedge clk) begin
	if (rs)
	Current_State <= S0;
	else
	Current_State <= Next_State;
end

always @(Current_State, t) begin
	case (Current_State)
	S0: Next_State = (t == 0) ? S1 : S0;
	S1: Next_State = (t == 0) ? S2 : S1;
	S2: Next_State = (t == 0) ? S3 : S2;
	S3: Next_State = (t == 0) ? S0 : S3;
	default: Next_State = S0;
	endcase
end

always @(posedge clk) begin
	if (rs) begin
		out_1 <= 3'b010;
		out_2 <= 3'b100;
	end else if (t == 0) begin
		case (Next_State)
		S0: begin out_1 <= 3'b010; out_2 <= 3'b100; end
		S1: begin out_1 <= 3'b001; out_2 <= 3'b100; end
		S2: begin out_1 <= 3'b100; out_2 <= 3'b010; end
		S3: begin out_1 <= 3'b100; out_2 <= 3'b001; end
		default: begin out_1 <= 3'b010; out_2 <= 3'b100; end
	endcase
	end
end

endmodule

