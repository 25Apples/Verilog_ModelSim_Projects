`timescale 1ns/1ps
module Nhat_testbench_D_FF_with_PRE_CLR();
reg PRE, CLR, CLK, D;
wire Q, Qn;

D_FF_with_PRE_CLR uut(
.PRE(PRE), .CLR(CLR), .CLK(CLK), .D(D),
.Q(Q), .Qn(Qn));

initial begin
	CLK = 0;
	PRE = 0;
	CLR = 0;
	D = 0;
end

always forever #5 CLK = ~CLK;
always forever #10 PRE = ~PRE;
always forever #20 CLR = ~CLR;
always forever #40 D = ~D;

endmodule
