module FullAdder (
input wire A, B, Cin, 
output wire S, Cout
);

assign S = A ^ B ^ Cin;
assign Cout = (A & B) | (Cin & ( A ^ B));

endmodule 

module RippleCarryAdder (
input wire [3:0] A, B, 
input wire Cin,
output wire [4:0] S
);

wire C1, C2, C3, Cout;
FullAdder FA0 (.A(A[0]), .B(B[0]), .Cin(Cin), .S(S[0]), .Cout(C1));
FullAdder FA1 (.A(A[1]), .B(B[1]), .Cin(C1), .S(S[1]), .Cout(C2));
FullAdder FA2 (.A(A[2]), .B(B[2]), .Cin(C2), .S(S[2]), .Cout(C3));
FullAdder FA3 (.A(A[3]), .B(B[3]), .Cin(C3), .S(S[3]), .Cout(Cout));
assign S[4] = Cout;

endmodule

